library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity hardware_FIFO is
  port (
    w_data: IN 
  
  );
end entity hardware_FIFO;



architecture beh of hardware_FIFO is
  component 

begin
  
      
  
end architecture beh;
